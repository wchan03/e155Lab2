// Wava Chan
// wchan@g.hmc.edu
// Sept. 4, 2025
// Top Level Module for Lab 2: Mutiplexed 7-Seg Display
// This module TODO: FINISH This

module lab2_wc(input logic clk, reset
                input logic [3:0] s1, s2, // Two DIP switches
                output logic [6:0] seg_disp1, seg_disp2);

                // Segment Display Module


                //TO DO 
                // Module (?) to drive the switching between two pins
                